-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 17.1.0 Build 590 10/25/2017 SJ Lite Edition
-- Created on Mon May 04 12:23:55 2020

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SeqDetFSM IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        Xin : IN STD_LOGIC := '0';
        Yout : OUT STD_LOGIC
    );
END SeqDetFSM;

ARCHITECTURE BEHAVIOR OF SeqDetFSM IS
    TYPE type_fstate IS (S0,S1,S2,S3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Xin)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= S0;
            Yout <= '0';
        ELSE
            Yout <= '0';
            CASE fstate IS
                WHEN S0 =>
                    IF ((Xin = '0')) THEN
                        reg_fstate <= S0;
                    ELSIF ((Xin = '1')) THEN
                        reg_fstate <= S1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S0;
                    END IF;

                    Yout <= '0';
                WHEN S1 =>
                    IF ((Xin = '0')) THEN
                        reg_fstate <= S2;
                    ELSIF ((Xin = '1')) THEN
                        reg_fstate <= S1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S1;
                    END IF;

                    Yout <= '0';
                WHEN S2 =>
                    IF ((Xin = '0')) THEN
                        reg_fstate <= S3;
                    ELSIF ((Xin = '1')) THEN
                        reg_fstate <= S1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S2;
                    END IF;

                    Yout <= '0';
                WHEN S3 =>
                    IF ((Xin = '0')) THEN
                        reg_fstate <= S0;
								Yout <= '0';
                    ELSIF ((Xin = '1')) THEN
                        reg_fstate <= S1;
								Yout <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S3;
                    END IF;
                WHEN OTHERS => 
                    Yout <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
